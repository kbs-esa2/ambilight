
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY framebuffer IS
PORT (

);
END framebuffer;

ARCHITECTURE framebuffer_rtl OF framebuffer IS



BEGIN

END MBlight_rtl;