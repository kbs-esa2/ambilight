
module PLL (
	clkin_clk,
	reset_reset,
	clkout_clk);	

	input		clkin_clk;
	input		reset_reset;
	output		clkout_clk;
endmodule
