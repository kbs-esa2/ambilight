// PLL.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module PLL (
		input  wire  clkin_clk,   //  clkin.clk
		output wire  clkout_clk,  // clkout.clk
		input  wire  reset_reset  //  reset.reset
	);

	PLL_altpll_0 altpll_0 (
		.clk                (clkin_clk),   //       inclk_interface.clk
		.reset              (reset_reset), // inclk_interface_reset.reset
		.read               (),            //             pll_slave.read
		.write              (),            //                      .write
		.address            (),            //                      .address
		.readdata           (),            //                      .readdata
		.writedata          (),            //                      .writedata
		.c0                 (clkout_clk),  //                    c0.clk
		.scandone           (),            //           (terminated)
		.scandataout        (),            //           (terminated)
		.areset             (1'b0),        //           (terminated)
		.locked             (),            //           (terminated)
		.phasedone          (),            //           (terminated)
		.phasecounterselect (4'b0000),     //           (terminated)
		.phaseupdown        (1'b0),        //           (terminated)
		.phasestep          (1'b0),        //           (terminated)
		.scanclk            (1'b0),        //           (terminated)
		.scanclkena         (1'b0),        //           (terminated)
		.scandata           (1'b0),        //           (terminated)
		.configupdate       (1'b0)         //           (terminated)
	);

endmodule
